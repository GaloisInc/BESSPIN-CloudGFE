package AWS_BSV_Top_Defs_Platform;

// ================================================================
// This package contains definitions of any platform-specific types
// and constants.

typedef 4  Num_DDR4;
typedef 2  Num_glcount;
typedef 16 Num_vDIP;
typedef 16 Num_vLED;

Bit #(64) ddr4_size = 'h_4_0000_0000; // 16 GB

// ================================================================

endpackage
