package AWS_BSV_Top_Defs_Platform;

// ================================================================
// This package contains definitions of any platform-specific types
// and constants.

typedef 2  Num_DDR4;
typedef 0  Num_glcount;
typedef 0  Num_vDIP;
typedef 0  Num_vLED;

Bit #(64) ddr4_size = 'h_8000_0000; // 2 GB

// ================================================================

endpackage
